module memory_ctrl #(
)(
)

endmodule
